// Instruction _ Mode definition

`define     MODE_IDLE   'd0
`define     MODE_SL     'd1
`define     MODE_RL     'd2
`define     MODE_WL     'd3
`define     MODE_PWM    'd4
`define     MODE_RS_ANI 8'b11000101
`define     MODE_RS_PIC 8'b10000101



// LED Color define

`define     COLOR_GREEN     3'b011
`define     COLOR_BLUE      3'b110
`define     COLOR_RED       3'b101
`define     COLOR_ORANGE    3'b001
`define     COLOR_OFF       3'b111


