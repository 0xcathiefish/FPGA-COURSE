// Version 1.0

`define ST_INS_IDLE         'd0
`define ST_INS_FETCH        'd1
`define ST_INS_ASSEMBLE     'd2
`define ST_INS_EXCUTE       'd3
`define ST_INS_DONE         'd4